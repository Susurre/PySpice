Modified Nodel Analysis Circuit
*Lecture 6 Circuit I
R1 1 2 5000k
R2 2 0 10
Vsrc 1 0 1
Isrc 0 2 1
.dc Vsrc 0 10 1
.ends