R+diode circuit to observe convergence of diode stamp
*from Lecture8 page43
v1 1 0 1 1 tran sin (1)
r1 1 2 1n
d1 2 0 somemodel
.tran 0.01 2 0
.end


