Modified Nodel Analysis Circuit
*Lecture 6 Circuit II Page-9
*if solver is V1=65.82V, V2=71.90V,
*then stamping for G is correct.
R1 1 0 5
G2 1 0 1 2 2
R3 1 2 6
R4 2 0 8
Is 0 2 10
*also, demo for .print command
.END