lc oscillation
c1 1 0 1 ic=1
l1 1 0 1
.tran 0.1 100 0.0
.end

